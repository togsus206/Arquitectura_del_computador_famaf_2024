`timescale 1ns / 1ps

module alu_tb();
	 parameter N = 64; // Ancho de datos de prueba
    logic clk;
    logic [N-1:0] a, b;
    logic [3:0] ALUControl;
    logic [N-1:0] result;
    logic zero_expected;

    // Instancia el módulo alu
    alu #(N) dut(a, b, ALUControl, result, zero);
		
    // Genera señal de reloj
    always begin
        clk = 0; #5; clk = 1; #5;
    end

    // Test de todas las operaciones
    initial begin
        $display("Test de todas las operaciones:");

        // Test de suma (positivo + positivo)
        a = 4'b0101;
        b = 4'b0010;
        ALUControl = 4'b0010;
        zero_expected = 0;
        #10;
        check_result("Suma (positivo + positivo)", zero_expected);

        // Test de resta (positivo - positivo)
        a = 4'b0101;
        b = 4'b0010;
        ALUControl = 4'b0110;
        zero_expected = 0;
        #10;
        check_result("Resta (positivo - positivo)", zero_expected);

        // Test de suma (negativo + negativo)
        a = 4'b1101;
        b = 4'b1010;
        ALUControl = 4'b0010;
        zero_expected = 0;
        #10;
        check_result("Suma (negativo + negativo)", zero_expected);

        // Test de resta (negativo - negativo)
        a = 4'b1101;
        b = 4'b1010;
        ALUControl = 4'b0110;
        zero_expected = 0;
        #10;
        check_result("Resta (negativo - negativo)", zero_expected);

        // Test de suma (positivo + negativo)
        a = 4'b0101;
        b = 4'b1010;
        ALUControl = 4'b0010;
        zero_expected = 1;
        #10;
        check_result("Suma (positivo + negativo)", zero_expected);

        // Test de resta (positivo - negativo)
        a = 4'b0101;
        b = 4'b1010;
        ALUControl = 4'b0110;
        zero_expected = 0;
        #10;
        check_result("Resta (positivo - negativo)", zero_expected);

        // Test de suma (negativo + positivo)
        a = 4'b1101;
        b = 4'b0010;
        ALUControl = 4'b0010;
        zero_expected = 0;
        #10;
        check_result("Suma (negativo + positivo)", zero_expected);

        // Test de resta (negativo - positivo)
        a = 4'b1101;
        b = 4'b0010;
        ALUControl = 4'b0110;
        zero_expected = 0;
        #10;
        check_result("Resta (negativo - positivo)", zero_expected);

        $finish;
    end

    // Función para verificar el resultado y la bandera zero
    function void check_result(string operation, logic zero_expected);
        if (result == 0 && zero_expected == 1)
            $display("%s: PASSED (Result = %h, Zero = %b)", operation, result, zero_expected);
        else if (result != 0 && zero_expected == 0)
            $display("%s: PASSED (Result = %h, Zero = %b)", operation, result, zero_expected);
        else
            $display("%s: FAILED (Result = %h, Zero = %b)", operation, result, zero_expected);
    endfunction

endmodule